/home/shadab/shadab/FPR/lef/all.lef